module project2-top (
);

endmodule
