module stopwatch (
);

endmodule
