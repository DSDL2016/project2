// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Thu May 19 17:04:13 2016

// synthesis message_off 10175

`timescale 1ns/1ns

module key_logic_fsm (
    clock,reset,k3,k1,
    run_timer,reset_timer);

    input clock;
    input reset;
    input k3;
    input k1;
    tri0 reset;
    tri0 k3;
    tri0 k1;
    output run_timer;
    output reset_timer;
    reg run_timer;
    reg reset_timer;
    reg [6:0] fstate;
    reg [6:0] reg_fstate;
    parameter s_pre_start=0,s_run=1,s_pre_pause=2,s_pause=3,s_idle=4,s_pre_reset=5,s_reset=6;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or k3 or k1)
    begin
        if (reset) begin
            reg_fstate <= s_idle;
            run_timer <= 1'b0;
            reset_timer <= 1'b0;
        end
        else begin
            run_timer <= 1'b0;
            reset_timer <= 1'b0;
            case (fstate)
                s_pre_start: begin
                    if ((~(k3) & ~(k1)))
                        reg_fstate <= s_run;
                    else if ((k3 & ~(k1)))
                        reg_fstate <= s_pre_start;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s_pre_start;

                    run_timer <= 1'b1;
                end
                s_run: begin
                    if ((k3 & ~(k1)))
                        reg_fstate <= s_pre_pause;
                    else if ((~(k3) & ~(k1)))
                        reg_fstate <= s_run;
                    else if ((~(k3) & k1))
                        reg_fstate <= s_pre_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s_run;

                    run_timer <= 1'b1;
                end
                s_pre_pause: begin
                    if ((~(k3) & ~(k1)))
                        reg_fstate <= s_pause;
                    else if ((k3 & ~(k1)))
                        reg_fstate <= s_pre_pause;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s_pre_pause;
                end
                s_pause: begin
                    if ((k3 & ~(k1)))
                        reg_fstate <= s_pre_start;
                    else if ((~(k3) & ~(k1)))
                        reg_fstate <= s_pause;
                    else if ((~(k3) & k1))
                        reg_fstate <= s_pre_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s_pause;
                end
                s_idle: begin
                    if ((k3 & ~(k1)))
                        reg_fstate <= s_pre_start;
                    else if ((~(k3) & ~(k1)))
                        reg_fstate <= s_idle;
                    else if ((~(k3) & k1))
                        reg_fstate <= s_pre_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s_idle;
                end
                s_pre_reset: begin
                    if ((~(k3) & k1))
                        reg_fstate <= s_pre_reset;
                    else if ((~(k3) & ~(k1)))
                        reg_fstate <= s_reset;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s_pre_reset;
                end
                s_reset: begin
                    reg_fstate <= s_idle;

                    reset_timer <= 1'b1;
                end
                default: begin
                    run_timer <= 1'bx;
                    reset_timer <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // key_logic_fsm
